-------------------------------------------------------------------------------
--
-- Title       : TanhL
-- Design      : TanhJoao
-- Author      : GCEM
-- Company     : nenhuma
--
-------------------------------------------------------------------------------
--
-- File        : TanhL.vhd
-- Generated   : Wed Apr 27 11:13:33 2016
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {TanhL} architecture {TanhL}}

library ieee;
use ieee.numeric_std.all;  
use IEEE.STD_LOGIC_1164.ALL;

entity TanhL is
	 port(
		 INPUT : in STD_LOGIC_VECTOR(24 downto 0);
		 OUTPUT : out STD_LOGIC_VECTOR(15 downto 0)
	     );
end TanhL;

--}} End of automatically maintained section

architecture TanhL of TanhL is	 

COMPONENT Func1Grau IS
	 port(
		 A      : in  STD_LOGIC_VECTOR(24 downto 0);
		 B      : in  STD_LOGIC_VECTOR(49 downto 0);
		 X      : in  STD_LOGIC_VECTOR(24 downto 0);
		 RESULT : out STD_LOGIC_VECTOR(15 downto 0));  
		 
END COMPONENT;	  

	SIGNAL AAux, XAux, TEMP1 : STD_LOGIC_VECTOR(24 DOWNTO 0); 
	SIGNAL BAux, TEMP0       : STD_LOGIC_VECTOR(49 DOWNTO 0); 
	SIGNAL SAIDAAux          : STD_LOGIC_VECTOR(15 DOWNTO 0); 		  
	SIGNAL OUTPUTAux0        : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL OUTPUTAux1        : STD_LOGIC_VECTOR(15 DOWNTO 0);          
begin 
	
	R0:	Func1Grau PORT MAP(A => AAux, B=> BAux, X=> XAux, RESULT=> SAIDAAux);	
	
	TEMP0 <= STD_LOGIC_VECTOR(SIGNED(INPUT) * "1111111110000000000000000");	   -- 'COMPLEMENTO DE DOIS'
	TEMP1 <= TEMP0(40) & TEMP0(39 DOWNTO 32) & TEMP0(31 DOWNTO 16);			   -- 'VALOR POSITIVO SE ENTRADA NEGATIVA'
	
	XAux <= INPUT WHEN INPUT(24) = '0' ELSE  
		    TEMP1 WHEN INPUT(24) = '1' ELSE	                                   -- VALOR JA COMPLEMENTADO   
			"0000000000000000000000000"; 

	BAux <= "00000000000000000000000000000000000000000000000000" WHEN XAux >= "0000000000000000000000000" AND  -- RETA 01
			XAux <= "0000000000111101100001000"	ELSE
		 
		    "00000000000000000000011001110110110000000000000000" WHEN XAUX >  "0000000000111101100001000" AND  -- RETA 02
			XAux <= "0000000001011001010010101"	ELSE
		 
		    "00000000000000000000111100100110000000000000000000" WHEN XAUX >  "0000000001011001010010101" AND  -- RETA 03
			XAux <= "0000000010000000000000000"	ELSE			
		 
		    "00000000000000000001101011000111000000000000000000" WHEN XAUX >  "0000000010000000000000000" AND  -- RETA 04
			XAux <= "0000000010100001110010101"	ELSE				
		 
		    "00000000000000000010010111001110000000000000000000" WHEN XAUX >  "0000000010100001110010101" AND  -- RETA 05
			XAux <= "0000000011001100110011001"	ELSE			
		 
		    "00000000000000000010111110001110110000000000000000" WHEN XAUX >  "0000000011001100110011001" AND  -- RETA 06
			XAux <= "0000000011111000010101010"	ELSE				
		 
		    "00000000000000000011011100010010010000000000000000" WHEN XAUX >  "0000000011111000010101010" AND  -- RETA 07
			XAux <= "0000000100110111100011010"	ELSE
		 
		    "00000000000000000011110000110100010000000000000000" WHEN XAUX >  "0000000100110111100011010" AND  -- RETA 08
			XAux <= "0000000110000000000000000"	ELSE					
		 
		    "00000000000000000011111100111001110000000000000000" WHEN XAUX >  "0000000110000000000000000" AND  -- RETA 09
			XAux <= "0000001010000000000000000"	ELSE	
			
			"00000000000000000000000000000000000000000000000000";
			
	AAux <= "0000000001110111000000111" WHEN XAux >= "0000000000000000000000000" AND  -- RETA 01
			XAux <= "0000000000111101100001000"	ELSE
		 
		    "0000000001011100000100100" WHEN XAUX >  "0000000000111101100001000" AND  -- RETA 02
			XAux <= "0000000001011001010010101"	ELSE
		 
		    "0000000001000011001011001" WHEN XAUX >  "0000000001011001010010101" AND  -- RETA 03
			XAux <= "0000000010000000000000000"	ELSE			
		 
		    "0000000000101011111010101" WHEN XAUX >  "0000000010000000000000000" AND  -- RETA 04
			XAux <= "0000000010100001110010101"	ELSE				
		 
		    "0000000000011010011110000" WHEN XAUX >  "0000000010100001110010101" AND  -- RETA 05
			XAux <= "0000000011001100110011001"	ELSE			
		 
		    "0000000000001110010000100" WHEN XAUX >  "0000000011001100110011001" AND  -- RETA 06
			XAux <= "0000000011111000010101010"	ELSE				
		 
		    "0000000000000110100001110" WHEN XAUX >  "0000000011111000010101010" AND  -- RETA 07
			XAux <= "0000000100110111100011010"	ELSE
		 
		    "0000000000000010010100010" WHEN XAUX >  "0000000100110111100011010" AND  -- RETA 08
			XAux <= "0000000110000000000000000"	ELSE					
		 
		    "0000000000000000010011101" WHEN XAUX >  "0000000110000000000000000" AND  -- RETA 09
			XAux <= "0000001010000000000000000"	ELSE	
			
			"0000000000000000000000000";	
	
	OUTPUTAux0 <=  STD_LOGIC_VECTOR(SIGNED(SAIDAAux) * "1110000000000000");	
	OUTPUTAux1 <=  OUTPUTAux0(31) &  OUTPUTAux0(27 DOWNTO 26) & OUTPUTAux0(25 DOWNTO 13); 
	
	OUTPUT <= SAIDAAux   WHEN INPUT(24) = '0' ELSE
			  OUTPUTAux1 WHEN INPUT(24) = '1' ELSE
			  "0000000000000000";	  
		  
end TanhL;
