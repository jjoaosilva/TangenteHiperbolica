-------------------------------------------------------------------------------
--
-- Title       : Somador
-- Design      : TanhJoao
-- Author      : GCEM
-- Company     : nenhuma
--
-------------------------------------------------------------------------------
--
-- File        : Somador.vhd
-- Generated   : Wed Apr 27 11:19:24 2016
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.20
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Somador} architecture {Somador}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Somador is
	 port(
		 INPUT1S : in STD_LOGIC_VECTOR(49 downto 0);
		 INPUT2S : in STD_LOGIC_VECTOR(49 downto 0);
		 RESULTS : out STD_LOGIC_VECTOR(50 downto 0)
	     );
end Somador;   

architecture Somador of Somador is 

COMPONENT HalfAdder IS
	 port(
		 INPUTA   : in STD_LOGIC;
		 INPUTB   : in STD_LOGIC;
		 CARRYIn  : in STD_LOGIC;
		 OUTPUT   : out STD_LOGIC;
		 CARRYOut : out STD_LOGIC);	 
END COMPONENT;

		SIGNAL TEMP: STD_LOGIC_VECTOR (49 downto 0) := "00000000000000000000000000000000000000000000000000";
		SIGNAL C   : STD_LOGIC_VECTOR (49 downto 0) := "00000000000000000000000000000000000000000000000000";

begin		   

HA0 : HALFADDER PORT MAP(INPUTA=> INPUT1S(0) , INPUTB=> INPUT2S(0) , CARRYIn=> '0'  , OUTPUT=> TEMP(0) , CARRYOut=> C(0) );
HA1 : HALFADDER PORT MAP(INPUTA=> INPUT1S(1) , INPUTB=> INPUT2S(1) , CARRYIn=> C(0) , OUTPUT=> TEMP(1) , CARRYOut=> C(1) );
HA2 : HALFADDER PORT MAP(INPUTA=> INPUT1S(2) , INPUTB=> INPUT2S(2) , CARRYIn=> C(1) , OUTPUT=> TEMP(2) , CARRYOut=> C(2) ); 
HA3 : HALFADDER PORT MAP(INPUTA=> INPUT1S(3) , INPUTB=> INPUT2S(3) , CARRYIn=> C(2) , OUTPUT=> TEMP(3) , CARRYOut=> C(3) ); 
HA4 : HALFADDER PORT MAP(INPUTA=> INPUT1S(4) , INPUTB=> INPUT2S(4) , CARRYIn=> C(3) , OUTPUT=> TEMP(4) , CARRYOut=> C(4) );
HA5 : HALFADDER PORT MAP(INPUTA=> INPUT1S(5) , INPUTB=> INPUT2S(5) , CARRYIn=> C(4) , OUTPUT=> TEMP(5) , CARRYOut=> C(5) );
HA6 : HALFADDER PORT MAP(INPUTA=> INPUT1S(6) , INPUTB=> INPUT2S(6) , CARRYIn=> C(5) , OUTPUT=> TEMP(6) , CARRYOut=> C(6) );
HA7 : HALFADDER PORT MAP(INPUTA=> INPUT1S(7) , INPUTB=> INPUT2S(7) , CARRYIn=> C(6) , OUTPUT=> TEMP(7) , CARRYOut=> C(7) );
HA8 : HALFADDER PORT MAP(INPUTA=> INPUT1S(8) , INPUTB=> INPUT2S(8) , CARRYIn=> C(7) , OUTPUT=> TEMP(8) , CARRYOut=> C(8) ); 
HA9 : HALFADDER PORT MAP(INPUTA=> INPUT1S(9) , INPUTB=> INPUT2S(9) , CARRYIn=> C(8) , OUTPUT=> TEMP(9) , CARRYOut=> C(9) ); 
HA10: HALFADDER PORT MAP(INPUTA=> INPUT1S(10), INPUTB=> INPUT2S(10), CARRYIn=> C(9) , OUTPUT=> TEMP(10), CARRYOut=> C(10)); 
HA11: HALFADDER PORT MAP(INPUTA=> INPUT1S(11), INPUTB=> INPUT2S(11), CARRYIn=> C(10), OUTPUT=> TEMP(11), CARRYOut=> C(11)); 
HA12: HALFADDER PORT MAP(INPUTA=> INPUT1S(12), INPUTB=> INPUT2S(12), CARRYIn=> C(11), OUTPUT=> TEMP(12), CARRYOut=> C(12)); 
HA13: HALFADDER PORT MAP(INPUTA=> INPUT1S(13), INPUTB=> INPUT2S(13), CARRYIn=> C(12), OUTPUT=> TEMP(13), CARRYOut=> C(13)); 
HA14: HALFADDER PORT MAP(INPUTA=> INPUT1S(14), INPUTB=> INPUT2S(14), CARRYIn=> C(13), OUTPUT=> TEMP(14), CARRYOut=> C(14)); 
HA15: HALFADDER PORT MAP(INPUTA=> INPUT1S(15), INPUTB=> INPUT2S(15), CARRYIn=> C(14), OUTPUT=> TEMP(15), CARRYOut=> C(15)); 
HA16: HALFADDER PORT MAP(INPUTA=> INPUT1S(16), INPUTB=> INPUT2S(16), CARRYIn=> C(15), OUTPUT=> TEMP(16), CARRYOut=> C(16));
HA17: HALFADDER PORT MAP(INPUTA=> INPUT1S(17), INPUTB=> INPUT2S(17), CARRYIn=> C(16), OUTPUT=> TEMP(17), CARRYOut=> C(17));
HA18: HALFADDER PORT MAP(INPUTA=> INPUT1S(18), INPUTB=> INPUT2S(18), CARRYIn=> C(17), OUTPUT=> TEMP(18), CARRYOut=> C(18));
HA19: HALFADDER PORT MAP(INPUTA=> INPUT1S(19), INPUTB=> INPUT2S(19), CARRYIn=> C(18), OUTPUT=> TEMP(19), CARRYOut=> C(19));
HA20: HALFADDER PORT MAP(INPUTA=> INPUT1S(20), INPUTB=> INPUT2S(20), CARRYIn=> C(19), OUTPUT=> TEMP(20), CARRYOut=> C(20));
HA21: HALFADDER PORT MAP(INPUTA=> INPUT1S(21), INPUTB=> INPUT2S(21), CARRYIn=> C(20), OUTPUT=> TEMP(21), CARRYOut=> C(21));
HA22: HALFADDER PORT MAP(INPUTA=> INPUT1S(22), INPUTB=> INPUT2S(22), CARRYIn=> C(21), OUTPUT=> TEMP(22), CARRYOut=> C(22));
HA23: HALFADDER PORT MAP(INPUTA=> INPUT1S(23), INPUTB=> INPUT2S(23), CARRYIn=> C(22), OUTPUT=> TEMP(23), CARRYOut=> C(23));
HA24: HALFADDER PORT MAP(INPUTA=> INPUT1S(24), INPUTB=> INPUT2S(24), CARRYIn=> C(23), OUTPUT=> TEMP(24), CARRYOut=> C(24));
HA25: HALFADDER PORT MAP(INPUTA=> INPUT1S(25), INPUTB=> INPUT2S(25), CARRYIn=> C(24), OUTPUT=> TEMP(25), CARRYOut=> C(25));
HA26: HALFADDER PORT MAP(INPUTA=> INPUT1S(26), INPUTB=> INPUT2S(26), CARRYIn=> C(25), OUTPUT=> TEMP(26), CARRYOut=> C(26));
HA27: HALFADDER PORT MAP(INPUTA=> INPUT1S(27), INPUTB=> INPUT2S(27), CARRYIn=> C(26), OUTPUT=> TEMP(27), CARRYOut=> C(27));
HA28: HALFADDER PORT MAP(INPUTA=> INPUT1S(28), INPUTB=> INPUT2S(28), CARRYIn=> C(27), OUTPUT=> TEMP(28), CARRYOut=> C(28));
HA29: HALFADDER PORT MAP(INPUTA=> INPUT1S(29), INPUTB=> INPUT2S(29), CARRYIn=> C(28), OUTPUT=> TEMP(29), CARRYOut=> C(29));
HA30: HALFADDER PORT MAP(INPUTA=> INPUT1S(30), INPUTB=> INPUT2S(30), CARRYIn=> C(29), OUTPUT=> TEMP(30), CARRYOut=> C(30));
HA31: HALFADDER PORT MAP(INPUTA=> INPUT1S(31), INPUTB=> INPUT2S(31), CARRYIn=> C(30), OUTPUT=> TEMP(31), CARRYOut=> C(31));
HA32: HALFADDER PORT MAP(INPUTA=> INPUT1S(32), INPUTB=> INPUT2S(32), CARRYIn=> C(31), OUTPUT=> TEMP(32), CARRYOut=> C(32));
HA33: HALFADDER PORT MAP(INPUTA=> INPUT1S(33), INPUTB=> INPUT2S(33), CARRYIn=> C(32), OUTPUT=> TEMP(33), CARRYOut=> C(33));
HA34: HALFADDER PORT MAP(INPUTA=> INPUT1S(34), INPUTB=> INPUT2S(34), CARRYIn=> C(33), OUTPUT=> TEMP(34), CARRYOut=> C(34));
HA35: HALFADDER PORT MAP(INPUTA=> INPUT1S(35), INPUTB=> INPUT2S(35), CARRYIn=> C(34), OUTPUT=> TEMP(35), CARRYOut=> C(35));
HA36: HALFADDER PORT MAP(INPUTA=> INPUT1S(36), INPUTB=> INPUT2S(36), CARRYIn=> C(35), OUTPUT=> TEMP(36), CARRYOut=> C(36));
HA37: HALFADDER PORT MAP(INPUTA=> INPUT1S(37), INPUTB=> INPUT2S(37), CARRYIn=> C(36), OUTPUT=> TEMP(37), CARRYOut=> C(37));
HA38: HALFADDER PORT MAP(INPUTA=> INPUT1S(38), INPUTB=> INPUT2S(38), CARRYIn=> C(37), OUTPUT=> TEMP(38), CARRYOut=> C(38));
HA39: HALFADDER PORT MAP(INPUTA=> INPUT1S(39), INPUTB=> INPUT2S(39), CARRYIn=> C(38), OUTPUT=> TEMP(39), CARRYOut=> C(39));
HA40: HALFADDER PORT MAP(INPUTA=> INPUT1S(40), INPUTB=> INPUT2S(40), CARRYIn=> C(39), OUTPUT=> TEMP(40), CARRYOut=> C(40));
HA41: HALFADDER PORT MAP(INPUTA=> INPUT1S(41), INPUTB=> INPUT2S(41), CARRYIn=> C(40), OUTPUT=> TEMP(41), CARRYOut=> C(41));
HA42: HALFADDER PORT MAP(INPUTA=> INPUT1S(42), INPUTB=> INPUT2S(42), CARRYIn=> C(41), OUTPUT=> TEMP(42), CARRYOut=> C(42));
HA43: HALFADDER PORT MAP(INPUTA=> INPUT1S(43), INPUTB=> INPUT2S(43), CARRYIn=> C(42), OUTPUT=> TEMP(43), CARRYOut=> C(43));
HA44: HALFADDER PORT MAP(INPUTA=> INPUT1S(44), INPUTB=> INPUT2S(44), CARRYIn=> C(43), OUTPUT=> TEMP(44), CARRYOut=> C(44));
HA45: HALFADDER PORT MAP(INPUTA=> INPUT1S(45), INPUTB=> INPUT2S(45), CARRYIn=> C(44), OUTPUT=> TEMP(45), CARRYOut=> C(45));
HA46: HALFADDER PORT MAP(INPUTA=> INPUT1S(46), INPUTB=> INPUT2S(46), CARRYIn=> C(45), OUTPUT=> TEMP(46), CARRYOut=> C(46));
HA47: HALFADDER PORT MAP(INPUTA=> INPUT1S(47), INPUTB=> INPUT2S(47), CARRYIn=> C(46), OUTPUT=> TEMP(47), CARRYOut=> C(47));
HA48: HALFADDER PORT MAP(INPUTA=> INPUT1S(48), INPUTB=> INPUT2S(48), CARRYIn=> C(47), OUTPUT=> TEMP(48), CARRYOut=> C(48));
HA49: HALFADDER PORT MAP(INPUTA=> INPUT1S(49), INPUTB=> INPUT2S(49), CARRYIn=> C(48), OUTPUT=> TEMP(49), CARRYOut=> C(49));	

	RESULTS <= C(49) & TEMP;

end Somador;
